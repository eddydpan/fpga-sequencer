module top (
    input logic clk,
    output logic LED,
    output logic RGB_R, 
    output logic RGB_G, 
    output logic RGB_B
);
    // top module


endmodule
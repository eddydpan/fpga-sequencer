`include "model.sv"
`include "button_matrix_controller.sv"
`include "audio_controller.sv"

module top(
    input logic clk,
    input logic _39a, 
    input logic _38b, 
    input logic _41a, 
    input logic _42b, // button col inputs
    output logic _36b, 
    output logic _37a, 
    output logic _29b, 
    output logic _31b, // row pin outputs for matrix scanning
    output logic _44b, // audio output pin
    output logic LED,
    output logic RGB_R, 
    output logic RGB_G, 
    output logic RGB_B
);
    localparam NUM_BEATS = 16;
    localparam BEATS_BUFFER = $clog2(NUM_BEATS)-1;
    // Instantiate model
    logic[6:0] data_in;
    logic[NUM_BEATS*4-1:0] beats; // 64 bit register: 16 beats x 4 bits each (pitch)
    logic[BEATS_BUFFER:0] beat_count; // 4 bits for 16 beats


    model #(
        .NUM_BEATS(NUM_BEATS)
    ) u_model (
        .clk(clk),
        .data_in(data_in),
        .beats(beats)
    );
    
    logic[3:0] button_index; // 4 bits for 16 buttons
    logic button_pressed;
    
    button_matrix_controller u_button_matrix_controller (
        .clk(clk),
        .col_inputs({_42b, _41a, _38b, _39a}),
        .row_outputs({_31b, _29b, _37a, _36b}),
        .button_index(button_index),
        .button_pressed(button_pressed)
    );

    audio_controller #(
        .NUM_BEATS(NUM_BEATS)
    ) u_audio_controller(
        .clk(clk),
        .beats(beats),
        .beat_count(beat_count),
        .pwm_out(_44b)
    );
    
    always_ff @(posedge clk) begin
        if (button_pressed) begin
            data_in <= {4'b0001, button_index}; // TODO: map pitch bits w/ rotary encoder #3
        end
        else begin
            // Cast modulo result to 4 bits (enough for values 0-8)
            data_in <= {BEATS_BUFFER'(beat_count % 9), beat_count};
        end
    end
    // Hardware debugger: Map button_index bits directly to LEDs
    // This will help debug what values are actually being detected
    always_comb begin
        if (button_pressed) begin
            // Map button_index bits to RGB and LED
            // bit[0] -> RGB_R (inverted: 0=on)
            // bit[1] -> RGB_G (inverted: 0=on)
            // bit[2] -> RGB_B (inverted: 0=on)
            // bit[3] -> LED (inverted: 0=on)
            RGB_R = ~button_index[0];
            RGB_G = ~button_index[1];
            RGB_B = ~button_index[2];
            LED = ~button_index[3];
        end else begin
            // No button pressed: all LEDs off (high)
            RGB_R = 1;
            RGB_G = 1;
            RGB_B = 1;
            LED = 1;
        end
    end

    

endmodule
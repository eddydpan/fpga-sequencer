`include "model.sv"
`include "button_matrix_controller.sv"
`include "audio_controller.sv"
`include "rotary_encoder.sv"
`include "seven_segment.sv"

module top(
    input logic clk,
    input logic _39a, 
    input logic _38b, 
    input logic _41a, 
    input logic _42b, // button col inputs
    output logic _36b, 
    output logic _37a, 
    output logic _29b, 
    output logic _31b, // row pin outputs for matrix scanning
    output logic _48b, // audio output pin
    //{_0a, _5a, _9b, _6a, _4a, _49a, _3b}
    output logic _9b, // seven segment display segments
    output logic _6a,
    output logic _4a,
    output logic _2a,
    output logic _0a,
    output logic _5a,
    output logic _3b,
    output logic _49a,
    input logic _45a, // rotary encoder button
    input logic _44b, // rotary encoder output B
    input logic _43a, // rotary encoder output A
    output logic LED,
    output logic RGB_R, 
    output logic RGB_G, 
    output logic RGB_B
);
    localparam PERIOD = 10'd4;
    localparam NUM_BEATS = 16;
    localparam BEATS_BUFFER = $clog2(NUM_BEATS);
    localparam CLK_FREQ = 12_000_000; // 12 MHz
    // Instantiate model
    logic [7:0] data_in;
    logic [NUM_BEATS*4-1:0] beats; // 64 bit register: 16 beats x 4 bits each (pitch)
    logic [BEATS_BUFFER-1:0] beat_count; // 4 bits for 16 beats
    logic [$clog2(CLK_FREQ)-1:0] clk_count = 0;
    logic [3:0] seconds;
    logic [3:0] note;

    logic [3:0] rotary_position;
    logic re_button_pressed;

    model #(
        .NUM_BEATS(NUM_BEATS)
    ) u_model (
        .clk(clk),
        .data_in(data_in),
        .beats(beats)
    );
    
    logic[3:0] button_index; // 4 bits for 16 buttons
    logic button_pressed;
    
    button_matrix_controller u_button_matrix_controller (
        .clk(clk),
        .col_inputs({_42b, _41a, _38b, _39a}),
        .row_outputs({_31b, _29b, _37a, _36b}),
        .button_index(button_index),
        .button_pressed(button_pressed)
    );

    rotary_encoder u_rotary_encoder(
        .clk(clk),
        .button(_45a),
        .signal_a(_43a),
        .signal_b(_44b),
        .button_pressed(re_button_pressed),
        .rotary_position(rotary_position)
    );

    audio_controller #(
        .CLK_FREQ(CLK_FREQ),
        .NUM_BEATS(NUM_BEATS),
        .PERIOD(PERIOD)
    ) u_audio_controller(
        .clk(clk),
        .beats(beats),
        .beat_count(beat_count),
        .pwm_out(_48b),
        .pitch (note)
    );

    seven_segment u_seven_segment (
        .clk(clk),
        .note (note),
        .seg_data({_0a, _5a, _9b, _6a, _4a, _49a, _3b}), // GFEDCBA
        .decimal(_2a)
    );
    
    always_ff @(posedge clk) begin
        // Increment seconds counter
        if (clk_count == CLK_FREQ - 1) begin
            seconds <= seconds + 1;
            clk_count <= 0;
        end else begin
            clk_count <= clk_count + 1;
        end

        if (button_pressed) begin
            // Concatenate rotary encoder position and button index to form data_in
            // data_in is {4 bits of pitch, 4 bits of beat index}
            data_in <= {rotary_position, button_index}; // TODO: map pitch bits w/ rotary encoder #3
        end

    end
    // Hardware debugger: Map button_index bits directly to LEDs
    // This will help debug what values are actually being detected
    always_comb begin
        if (button_pressed) begin
            // Map button_index bits to RGB and LED
            // bit[0] -> RGB_R (inverted: 0=on)
            // bit[1] -> RGB_G (inverted: 0=on)
            // bit[2] -> RGB_B (inverted: 0=on)
            // bit[3] -> LED (inverted: 0=on)
            RGB_R = ~button_index[0];
            RGB_G = ~button_index[1];
            RGB_B = ~button_index[2];
            LED = ~button_index[3];
        end else begin
            // No button pressed: all LEDs off (high)
            RGB_R = 1;
            RGB_G = 1;
            RGB_B = 1;
            LED = 1;
        end
    end

    

endmodule